module top_module( 
    input a, 
    input b, 
    output out );
    xnor x1(out,a,b);
endmodule
