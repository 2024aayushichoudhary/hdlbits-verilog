module xor_gate(
  input a,b,
  output out
);
  xor x1(out,a,b);
endmodule
