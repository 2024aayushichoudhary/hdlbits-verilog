// HDLBits: AND gate
// Topic: Basic Gates
module top_module( 
    input a, 
    input b, 
    output out );
    //and a1(out,a,b);
  assign out=a&b;

endmodule
